library verilog;
use verilog.vl_types.all;
entity final_counter_vlg_check_tst is
    port(
        tick            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end final_counter_vlg_check_tst;
