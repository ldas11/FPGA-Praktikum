library verilog;
use verilog.vl_types.all;
entity final_counter_vlg_vec_tst is
end final_counter_vlg_vec_tst;
